// Memory initialization for simulation
// Generated from machine code

0A 00 08 20 14 00 09 20 05 00 0A 20 20 58 09 01
22 60 6A 01
