// Memory initialization for simulation
// Generated from machine code

0A 00 08 20 14 00 09 20 05 00 0A 20 20 58 09 01
22 60 6A 01 03 00 28 11 64 00 0D 20 02 00 08 11
C8 00 0E 20 2C 01 0F 20 90 01 18 20
