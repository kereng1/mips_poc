2008000A  # ADDI $t0, $zero, 10      # $t0 = 10
20090014  # ADDI $t1, $zero, 20      # $t1 = 20
200A0005  # ADDI $t2, $zero, 5       # $t2 = 5
01095820  # ADD $t3, $t0, $t1        # $t3 = $t0 + $t1 = 10 + 20 = 30
016A6022  # SUB $t4, $t3, $t2        # $t4 = $t3 - $t2 = 30 - 5 = 25
